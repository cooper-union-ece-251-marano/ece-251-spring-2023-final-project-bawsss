///////////////////////////////////////////////////////////////////////////////
//
// ALU module header
//
// An alu module header for your Computer Architecture Elements Catalog
//
// module: alu
// hdl: Verilog
//
// author: Fred Kim <fred.kim@cooper.edu>
//
///////////////////////////////////////////////////////////////////////////////

`ifndef ALU_SVH
`define ALU_SVH

`define ALU_CTRL_AND 3'b000
`define ALU_CTRL_OR  3'b001
`define ALU_CTRL_ADD 3'b010
`define ALU_CTRL_SLL 3'b011
`define ALU_CTRL_NOR 3'b100
`define ALU_CTRL_SRL 3'b101
`define ALU_CTRL_SUB 3'b110
`define ALU_CTRL_SLT 3'b111

`endif // ALU_SVH
